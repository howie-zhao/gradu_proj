module tb_overall (
    
);

endmodule //tb_overall